`timescale 1 ns/100 ps
// Version: v12.4 12.900.0.16
// File used only for Simulation


module sdf_IOPAD_TRI(
       PAD,
       D,
       E
    );
output PAD;
input  D;
input  E;

    wire NET_OIN_VDD, NET_EIN_VDD;
    
    IOPAD_TRI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD)
        , .PAD_P(PAD));
    IOPAD_VDD U_VCCA (.OIN_P(D), .EIN_P(E), .IOUT_VDD(), .OIN_VDD(
        NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN());
    
endmodule


module sdf_IOPAD_IN(
       PAD,
       Y
    );
input  PAD;
output Y;

    wire NET_IOUT_VDD, NET_IOUT_IN, ADLIB_GND;
    wire GND_power_net1;
    assign ADLIB_GND = GND_power_net1;
    
    IOPAD_IN_VDDI U_VCCI (.PAD_P(PAD), .IOUT_VDD(NET_IOUT_VDD));
    IOPAD_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .IOUT_P(Y));
    IOPAD_VDD U_VCCA (.OIN_P(ADLIB_GND), .EIN_P(ADLIB_GND), .IOUT_VDD(
        NET_IOUT_VDD), .OIN_VDD(), .EIN_VDD(), .IOUT_IN(NET_IOUT_IN));
    GND GND_power_inst1 (.Y(GND_power_net1));
    
endmodule


module sdf_IOPAD_BI(
       PAD,
       D,
       E,
       Y
    );
inout  PAD;
input  D;
input  E;
output Y;

    wire NET_IOUT_VDD, NET_IOUT_IN, NET_OIN_VDD, NET_EIN_VDD;
    
    IOPAD_BI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), 
        .IOUT_VDD(NET_IOUT_VDD), .PAD_P(PAD));
    IOPAD_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .IOUT_P(Y));
    IOPAD_VDD U_VCCA (.OIN_P(D), .EIN_P(E), .IOUT_VDD(NET_IOUT_VDD), 
        .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN(
        NET_IOUT_IN));
    
endmodule


module demo_sb(
       DEVRST_N,
       GPIO_9_F2M,
       MMUART_0_RXD_F2M,
       SPI_0_DI,
       GPIO_2_M2F,
       GPIO_3_M2F,
       GPIO_4_M2F,
       GPIO_8_M2F,
       MMUART_0_TXD_M2F,
       SPI_0_DO,
       I2C_0_SCL,
       I2C_0_SDA,
       SPI_0_CLK,
       SPI_0_SS0
    );
input  DEVRST_N;
input  GPIO_9_F2M;
input  MMUART_0_RXD_F2M;
input  SPI_0_DI;
output GPIO_2_M2F;
output GPIO_3_M2F;
output GPIO_4_M2F;
output GPIO_8_M2F;
output MMUART_0_TXD_M2F;
output SPI_0_DO;
inout  I2C_0_SCL;
inout  I2C_0_SDA;
inout  SPI_0_CLK;
inout  SPI_0_SS0;

    wire BIBUF_0_Y, demo_sb_sb_0_I2C_0_SDA_M2F, BIBUF_1_Y, 
        demo_sb_sb_0_I2C_0_SCL_M2F, GPIO_9_F2M_c, MMUART_0_RXD_F2M_c, 
        GPIO_2_M2F_c, GPIO_3_M2F_c, GPIO_4_M2F_c, GPIO_8_M2F_c, 
        MMUART_0_TXD_M2F_c, demo_sb_sb_0_I2C_0_SDA_M2F_OE, 
        demo_sb_sb_0_I2C_0_SCL_M2F_OE, \demo_sb_sb_0/SYSRESET_POR_Z , 
        \demo_sb_sb_0/FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC , 
        \demo_sb_sb_0/LOCK , \demo_sb_sb_0/CORERESETP_0_RESET_N_F2M , 
        \demo_sb_sb_0/CORERESETP_0/POWER_ON_RESET_N_clk_base_Z , VCC, 
        \demo_sb_sb_0/CORERESETP_0/sm1_areset_n_q1_Z , GND, 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD_Y , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD_Y , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD_Y , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE , 
        \demo_sb_sb_0/CCC_0/GL0_net , ff_to_start_net, 
        \GPIO_3_M2F_obuf/U0/DOUT1 , \GPIO_3_M2F_obuf/U0/DOUT , 
        \GPIO_3_M2F_obuf/U0/EOUT1 , \GPIO_3_M2F_obuf/U0/EOUT , 
        \BIBUF_1/U0/DOUT1 , \BIBUF_1/U0/DOUT , \BIBUF_1/U0/EOUT1 , 
        \BIBUF_1/U0/EOUT , \BIBUF_1/U0/YIN1 , \BIBUF_1/U0/YIN , 
        \MMUART_0_RXD_F2M_ibuf/U0/YIN1 , 
        \MMUART_0_RXD_F2M_ibuf/U0/YIN , 
        \demo_sb_sb_0/CCC_0/CCC_INST/CLK0_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/CLK1_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/CLK2_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/CLK3_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX0_SEL_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX1_SEL_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX2_SEL_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX3_SEL_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX0_HOLD_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX1_HOLD_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX2_HOLD_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX3_HOLD_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX0_ARST_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX1_ARST_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX2_ARST_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX3_ARST_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PLL_BYPASS_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PLL_ARST_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PLL_POWERDOWN_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/GPD0_ARST_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/GPD1_ARST_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/GPD2_ARST_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/GPD3_ARST_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PRESET_N_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PCLK_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PSEL_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PENABLE_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWRITE_net , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[7] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[6] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[5] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[4] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[3] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[2] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[7] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[6] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[5] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[4] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[3] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[2] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[1] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/COLF_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CRSF_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2HCALIB_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDIF_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_DVF_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_ERRF_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_EV_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CLK_BASE_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_BREADY_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_RREADY_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WLAST_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WVALID_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PRESET_N_net , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD/YIN , 
        \MMUART_0_TXD_M2F_obuf/U0/DOUT1 , 
        \MMUART_0_TXD_M2F_obuf/U0/DOUT , 
        \MMUART_0_TXD_M2F_obuf/U0/EOUT1 , 
        \MMUART_0_TXD_M2F_obuf/U0/EOUT , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD/YIN , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD/YIN , 
        \GPIO_4_M2F_obuf/U0/DOUT1 , \GPIO_4_M2F_obuf/U0/DOUT , 
        \GPIO_4_M2F_obuf/U0/EOUT1 , \GPIO_4_M2F_obuf/U0/EOUT , 
        \GPIO_2_M2F_obuf/U0/DOUT1 , \GPIO_2_M2F_obuf/U0/DOUT , 
        \GPIO_2_M2F_obuf/U0/EOUT1 , \GPIO_2_M2F_obuf/U0/EOUT , 
        \GPIO_9_F2M_ibuf/U0/YIN1 , \GPIO_9_F2M_ibuf/U0/YIN , 
        \BIBUF_0/U0/DOUT1 , \BIBUF_0/U0/DOUT , \BIBUF_0/U0/EOUT1 , 
        \BIBUF_0/U0/EOUT , \BIBUF_0/U0/YIN1 , \BIBUF_0/U0/YIN , 
        \GPIO_8_M2F_obuf/U0/DOUT1 , \GPIO_8_M2F_obuf/U0/DOUT , 
        \GPIO_8_M2F_obuf/U0/EOUT1 , \GPIO_8_M2F_obuf/U0/EOUT , 
        \demo_sb_sb_0/SYSRESET_POR/UTDO_net , 
        \demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1_YR , 
        \demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1 , 
        \demo_sb_sb_0/CCC_0/GL0_INST/U0_YWn_GEast , AFLSDF_VCC, 
        AFLSDF_GND, AFLSDF_INV_0_net_1;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign AFLSDF_GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign AFLSDF_VCC = VCC_power_net1;
    
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_78  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_171  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_113  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_174  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_86  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[2] ), 
        .IPC());
    IOOUTFF_BYPASS \GPIO_4_M2F_obuf/U0/U_IOOUTFF  (.A(
        \GPIO_4_M2F_obuf/U0/DOUT1 ), .Y(\GPIO_4_M2F_obuf/U0/DOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_271  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_80  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_223  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_129  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_21  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_121  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net ), 
        .IPB(), .IPC());
    sdf_IOPAD_TRI \GPIO_3_M2F_obuf/U0/U_IOPAD  (.PAD(GPIO_3_M2F), .D(
        \GPIO_3_M2F_obuf/U0/DOUT ), .E(\GPIO_3_M2F_obuf/U0/EOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_170  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net )
        , .IPB(), .IPC());
    IOOUTFF_BYPASS \MMUART_0_TXD_M2F_obuf/U0/U_IOOUTFF  (.A(
        \MMUART_0_TXD_M2F_obuf/U0/DOUT1 ), .Y(
        \MMUART_0_TXD_M2F_obuf/U0/DOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_232  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_165  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_124  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_242  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_105  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[5] ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_221  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] )
        , .IPC());
    sdf_IOPAD_TRI \MMUART_0_TXD_M2F_obuf/U0/U_IOPAD  (.PAD(
        MMUART_0_TXD_M2F), .D(\MMUART_0_TXD_M2F_obuf/U0/DOUT ), .E(
        \MMUART_0_TXD_M2F_obuf/U0/EOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_167  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_234  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] )
        , .IPC());
    IOINFF_BYPASS 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD/U_IOINFF  (.A(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD_Y ), .Y(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD/YIN ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_112  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_107  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_244  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] ), 
        .IPC());
    SYSRESET_FF \demo_sb_sb_0/SYSRESET_POR/INST_SYSRESET_FF_IP  (
        .UDRCAP(), .UDRSH(), .UDRUPD(), .UIREG({nc0, nc1, nc2, nc3, 
        nc4, nc5, nc6, nc7}), .URSTB(), .UDRCK(), .UTDI(), 
        .POWER_ON_RESET_N(\demo_sb_sb_0/SYSRESET_POR_Z ), .FF_TO_START(
        ff_to_start_net), .FF_DONE(), .UTDO(
        \demo_sb_sb_0/SYSRESET_POR/UTDO_net ), .DEVRST_N(DEVRST_N), 
        .TDI(VCC), .TMS(VCC), .TCK(VCC), .TRSTB(VCC), .TDO());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_120  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_235  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_245  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_93  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_DVF_net ), 
        .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_53  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_14  (.A(VCC)
        , .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX2_ARST_N_net ), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/GPD0_ARST_N_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[4] ));
    CCC #( .INIT(210'h0000007FB8000044D74000307C6318C6318C61EC0404040400301)
        , .VCOFREQUENCY(800.000000) )  
        \demo_sb_sb_0/CCC_0/CCC_INST/INST_CCC_IP  (.Y0(), .Y1(), .Y2(), 
        .Y3(), .PRDATA({nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15}), 
        .LOCK(\demo_sb_sb_0/LOCK ), .BUSY(), .CLK0(
        \demo_sb_sb_0/CCC_0/CCC_INST/CLK0_net ), .CLK1(
        \demo_sb_sb_0/CCC_0/CCC_INST/CLK1_net ), .CLK2(
        \demo_sb_sb_0/CCC_0/CCC_INST/CLK2_net ), .CLK3(
        \demo_sb_sb_0/CCC_0/CCC_INST/CLK3_net ), .NGMUX0_SEL(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX0_SEL_net ), .NGMUX1_SEL(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX1_SEL_net ), .NGMUX2_SEL(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX2_SEL_net ), .NGMUX3_SEL(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX3_SEL_net ), .NGMUX0_HOLD_N(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX0_HOLD_N_net ), 
        .NGMUX1_HOLD_N(\demo_sb_sb_0/CCC_0/CCC_INST/NGMUX1_HOLD_N_net )
        , .NGMUX2_HOLD_N(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX2_HOLD_N_net ), 
        .NGMUX3_HOLD_N(\demo_sb_sb_0/CCC_0/CCC_INST/NGMUX3_HOLD_N_net )
        , .NGMUX0_ARST_N(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX0_ARST_N_net ), 
        .NGMUX1_ARST_N(\demo_sb_sb_0/CCC_0/CCC_INST/NGMUX1_ARST_N_net )
        , .NGMUX2_ARST_N(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX2_ARST_N_net ), 
        .NGMUX3_ARST_N(\demo_sb_sb_0/CCC_0/CCC_INST/NGMUX3_ARST_N_net )
        , .PLL_BYPASS_N(\demo_sb_sb_0/CCC_0/CCC_INST/PLL_BYPASS_N_net )
        , .PLL_ARST_N(\demo_sb_sb_0/CCC_0/CCC_INST/PLL_ARST_N_net ), 
        .PLL_POWERDOWN_N(
        \demo_sb_sb_0/CCC_0/CCC_INST/PLL_POWERDOWN_N_net ), 
        .GPD0_ARST_N(\demo_sb_sb_0/CCC_0/CCC_INST/GPD0_ARST_N_net ), 
        .GPD1_ARST_N(\demo_sb_sb_0/CCC_0/CCC_INST/GPD1_ARST_N_net ), 
        .GPD2_ARST_N(\demo_sb_sb_0/CCC_0/CCC_INST/GPD2_ARST_N_net ), 
        .GPD3_ARST_N(\demo_sb_sb_0/CCC_0/CCC_INST/GPD3_ARST_N_net ), 
        .PRESET_N(\demo_sb_sb_0/CCC_0/CCC_INST/PRESET_N_net ), .PCLK(
        \demo_sb_sb_0/CCC_0/CCC_INST/PCLK_net ), .PSEL(
        \demo_sb_sb_0/CCC_0/CCC_INST/PSEL_net ), .PENABLE(
        \demo_sb_sb_0/CCC_0/CCC_INST/PENABLE_net ), .PWRITE(
        \demo_sb_sb_0/CCC_0/CCC_INST/PWRITE_net ), .PADDR({
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[7] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[6] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[5] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[4] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[3] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[2] }), .PWDATA({
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[7] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[6] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[5] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[4] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[3] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[2] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[1] , 
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[0] }), .CLK0_PAD(GND), 
        .CLK1_PAD(GND), .CLK2_PAD(GND), .CLK3_PAD(GND), .GL0(), .GL1(), 
        .GL2(), .GL3(\demo_sb_sb_0/CCC_0/GL0_net ), .RCOSC_25_50MHZ(
        \demo_sb_sb_0/FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC )
        , .RCOSC_1MHZ(GND), .XTLOSC(GND));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_54  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_9  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/CCC_0/CCC_INST/PLL_BYPASS_N_net ), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX3_SEL_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[7] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_213  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_119  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_87  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[3] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_1  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net ), 
        .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_3  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_111  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] )
        , .IPC());
    IOENFF_BYPASS \GPIO_2_M2F_obuf/U0/U_IOENFF  (.A(
        \GPIO_2_M2F_obuf/U0/EOUT1 ), .Y(\GPIO_2_M2F_obuf/U0/EOUT ));
    sdf_IOPAD_IN \MMUART_0_RXD_F2M_ibuf/U0/U_IOPAD  (.PAD(
        MMUART_0_RXD_F2M), .Y(\MMUART_0_RXD_F2M_ibuf/U0/YIN1 ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_268  
        (.A(VCC), .B(\demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1_YR ), .C(VCC)
        , .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CLK_BASE_net ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_114  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_208  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_0  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_211  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_175  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_82  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] )
        , .IPC());
    SLE \demo_sb_sb_0/CORERESETP_0/sm1_areset_n_q1  (.D(VCC), .CLK(
        \demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1 ), .EN(
        VCC), .ALn(\demo_sb_sb_0/SYSRESET_POR_Z ), .ADn(VCC), .SLn(VCC)
        , .SD(GND), .LAT(GND), .Q(
        \demo_sb_sb_0/CORERESETP_0/sm1_areset_n_q1_Z ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_2  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_110  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_177  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_256  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_260  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_200  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_125  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_2  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(\demo_sb_sb_0/CCC_0/CCC_INST/PCLK_net ), 
        .IPB(\demo_sb_sb_0/CCC_0/CCC_INST/NGMUX0_SEL_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[0] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_127  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_65  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net )
        , .IPC());
    sdf_IOPAD_TRI \GPIO_2_M2F_obuf/U0/U_IOPAD  (.PAD(GPIO_2_M2F), .D(
        \GPIO_2_M2F_obuf/U0/DOUT ), .E(\GPIO_2_M2F_obuf/U0/EOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_286  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_43  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_44  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_156  
        (.A(GPIO_9_F2M_c), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_69  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] )
        , .IPC());
    INV_BA AFLSDF_INV_0 (.A(\demo_sb_sb_0/CCC_0/GL0_net ), .Y(
        AFLSDF_INV_0_net_1));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_73  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_278  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_81  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_74  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] )
        , .IPB(), .IPC());
    IOENFF_BYPASS \GPIO_4_M2F_obuf/U0/U_IOENFF  (.A(
        \GPIO_4_M2F_obuf/U0/EOUT1 ), .Y(\GPIO_4_M2F_obuf/U0/EOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_68  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_262  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_196  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] )
        , .IPC());
    IOINFF_BYPASS 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD/U_IOINFF  (.A(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD_Y ), .Y(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD/YIN ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_202  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/SYSRESET_POR/IP_INTERFACE_0  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\demo_sb_sb_0/SYSRESET_POR/UTDO_net ), 
        .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_264  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_228  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_186  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_115  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_1  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\demo_sb_sb_0/CCC_0/CCC_INST/CLK1_net ), 
        .IPB(\demo_sb_sb_0/CCC_0/CCC_INST/PENABLE_net ), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_204  
        (.A(VCC), .B(GND), .C(GND), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_270  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_RREADY_net ), 
        .IPC());
    IOIN_IB \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD/U_IOIN  (.YIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD/YIN ), .E(GND), .Y(
        ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_117  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] )
        , .IPC());
    sdf_IOPAD_IN \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD/U_IOPAD  
        (.PAD(SPI_0_DI), .Y(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD_Y ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_265  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_205  
        (.A(VCC), .B(GND), .C(GND), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WLAST_net ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_96  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CRSF_net ), .IPB(
        ), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_56  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_220  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_4  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX0_HOLD_N_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[2] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_90  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[6] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_50  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] )
        , .IPB(), .IPC());
    sdf_IOPAD_TRI \GPIO_8_M2F_obuf/U0/U_IOPAD  (.PAD(GPIO_8_M2F), .D(
        \GPIO_8_M2F_obuf/U0/DOUT ), .E(\GPIO_8_M2F_obuf/U0/EOUT ));
    IOINFF_BYPASS \BIBUF_0/U0/U_IOINFF  (.A(\BIBUF_0/U0/YIN1 ), .Y(
        \BIBUF_0/U0/YIN ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_158  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net )
        , .IPB(), .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_5  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX1_HOLD_N_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[3] ));
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_16  (.A(VCC)
        , .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/GPD2_ARST_N_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[6] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_257  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_0  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\demo_sb_sb_0/CCC_0/CCC_INST/CLK0_net ), 
        .IPB(\demo_sb_sb_0/CCC_0/CCC_INST/PSEL_net ), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_259  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_272  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_218  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_198  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_8  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_274  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_15  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_35  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_188  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_153  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_287  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_222  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_275  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PRESET_N_net ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_210  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_19  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_39  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] )
        , .IPC());
    sdf_IOPAD_BI \BIBUF_1/U0/U_IOPAD  (.PAD(I2C_0_SCL), .D(
        \BIBUF_1/U0/DOUT ), .E(\BIBUF_1/U0/EOUT ), .Y(
        \BIBUF_1/U0/YIN1 ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_224  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_193  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_25  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_97  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/COLF_net ), .IPB(
        ), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_57  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_18  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_38  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_46  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_225  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_183  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_40  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_29  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_152  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net )
        , .IPC());
    RGB_NG \demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1  (.An(
        \demo_sb_sb_0/CCC_0/GL0_INST/U0_YWn_GEast ), .ENn(GND), .YL(), 
        .YR(\demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1_YR ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_76  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] )
        , .IPC());
    IOINFF_BYPASS \BIBUF_1/U0/U_IOINFF  (.A(\BIBUF_1/U0/YIN1 ), .Y(
        \BIBUF_1/U0/YIN ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_236  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_92  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_ERRF_net ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_70  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_52  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_246  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_28  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_15  (.A(VCC)
        , .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX3_ARST_N_net ), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/GPD1_ARST_N_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[5] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_192  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_212  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_63  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] )
        , .IPC());
    RCOSC_25_50MHZ #( .FREQUENCY(50.000000) )  
        \demo_sb_sb_0/FABOSC_0/I_RCOSC_25_50MHZ  (.CLKOUT(
        \demo_sb_sb_0/FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_64  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_182  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_253  
        (.A(VCC), .B(VCC), .C(GND), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_214  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_159  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net )
        , .IPC());
    IOINFF_BYPASS \GPIO_9_F2M_ibuf/U0/U_IOINFF  (.A(
        \GPIO_9_F2M_ibuf/U0/YIN1 ), .Y(\GPIO_9_F2M_ibuf/U0/YIN ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_151  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_136  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_146  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_154  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_251  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_215  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_199  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] )
        , .IPC());
    IOOUTFF_BYPASS \GPIO_2_M2F_obuf/U0/U_IOOUTFF  (.A(
        \GPIO_2_M2F_obuf/U0/DOUT1 ), .Y(\GPIO_2_M2F_obuf/U0/DOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_47  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_283  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_91  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[7] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_51  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_194  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_150  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_189  
        (.A(BIBUF_0_Y), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_181  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_77  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_184  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_281  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] )
        , .IPC());
    IOOUTFF_BYPASS \BIBUF_1/U0/U_IOOUTFF  (.A(\BIBUF_1/U0/DOUT1 ), .Y(
        \BIBUF_1/U0/DOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_42  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_72  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_180  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net )
        , .IPB(), .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_11  (.A(VCC)
        , .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/CCC_0/CCC_INST/PLL_POWERDOWN_N_net ), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX3_HOLD_N_net ), .IPC());
    sdf_IOPAD_IN \GPIO_9_F2M_ibuf/U0/U_IOPAD  (.PAD(GPIO_9_F2M), .Y(
        \GPIO_9_F2M_ibuf/U0/YIN1 ));
    IP_INTERFACE ip_interface_inst (.A(VCC), .B(ff_to_start_net), .C(
        VCC), .IPA(), .IPB(), .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_3  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/CCC_0/CCC_INST/PRESET_N_net ), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX1_SEL_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[1] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_138  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_148  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net )
        , .IPC());
    sdf_IOPAD_BI \BIBUF_0/U0/U_IOPAD  (.PAD(I2C_0_SDA), .D(
        \BIBUF_0/U0/DOUT ), .E(\BIBUF_0/U0/EOUT ), .Y(
        \BIBUF_0/U0/YIN1 ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_85  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[1] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_237  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] )
        , .IPC());
    sdf_IOPAD_BI \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD/U_IOPAD  
        (.PAD(SPI_0_SS0), .D(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT )
        , .E(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE )
        , .Y(\demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD_Y ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_247  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_239  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_249  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] )
        , .IPC());
    IOINFF_BYPASS \MMUART_0_RXD_F2M_ibuf/U0/U_IOINFF  (.A(
        \MMUART_0_RXD_F2M_ibuf/U0/YIN1 ), .Y(
        \MMUART_0_RXD_F2M_ibuf/U0/YIN ));
    IOINFF_BYPASS 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD/U_IOINFF  (.A(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD_Y ), .Y(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD/YIN ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_89  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[5] ), 
        .IPC());
    IOIN_IB \GPIO_9_F2M_ibuf/U0/U_IOIN  (.YIN(\GPIO_9_F2M_ibuf/U0/YIN )
        , .E(GND), .Y(GPIO_9_F2M_c));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_155  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_13  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_41  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_33  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_266  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_14  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_34  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_206  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_9  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_5  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_157  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_133  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_88  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[4] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_143  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_71  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_195  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] )
        , .IPC());
    IOENFF_BYPASS \BIBUF_0/U0/U_IOENFF  (.A(\BIBUF_0/U0/EOUT1 ), .Y(
        \BIBUF_0/U0/EOUT ));
    IOIN_IB \MMUART_0_RXD_F2M_ibuf/U0/U_IOIN  (.YIN(
        \MMUART_0_RXD_F2M_ibuf/U0/YIN ), .E(GND), .Y(
        MMUART_0_RXD_F2M_c));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_66  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_197  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_23  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_60  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_185  
        (.A(MMUART_0_RXD_F2M_c), .B(BIBUF_1_Y), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_24  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_187  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_166  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_106  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_132  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_142  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net )
        , .IPC());
    IOENFF_BYPASS \MMUART_0_TXD_M2F_obuf/U0/U_IOENFF  (.A(
        \MMUART_0_TXD_M2F_obuf/U0/EOUT1 ), .Y(
        \MMUART_0_TXD_M2F_obuf/U0/EOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_258  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_276  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_233  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_243  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_139  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_250  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_4  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_149  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_131  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_141  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2HCALIB_net ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_134  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net ), 
        .IPB(), .IPC());
    IOENFF_BYPASS \BIBUF_1/U0/U_IOENFF  (.A(\BIBUF_1/U0/EOUT1 ), .Y(
        \BIBUF_1/U0/EOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_67  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_231  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_226  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_144  
        (.A(\demo_sb_sb_0/LOCK ), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net )
        , .IPB(), .IPC());
    IOTRI_OB_EB \GPIO_3_M2F_obuf/U0/U_IOTRI  (.D(GPIO_3_M2F_c), .E(VCC)
        , .DOUT(\GPIO_3_M2F_obuf/U0/DOUT1 ), .EOUT(
        \GPIO_3_M2F_obuf/U0/EOUT1 ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_7  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_8  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/CCC_0/CCC_INST/PWRITE_net ), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX2_SEL_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[6] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_241  
        (.A(VCC), .B(GND), .C(GND), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] ), 
        .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_BREADY_net ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_176  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_168  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_130  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_280  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_140  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_EV_net ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_108  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_62  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_267  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_17  (.A(VCC)
        , .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/GPD3_ARST_N_net ), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[7] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_269  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_207  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_13  (.A(VCC)
        , .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX1_ARST_N_net ), .IPB(), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[3] ));
    sdf_IOPAD_TRI \GPIO_4_M2F_obuf/U0/U_IOPAD  (.PAD(GPIO_4_M2F), .D(
        \GPIO_4_M2F_obuf/U0/DOUT ), .E(\GPIO_4_M2F_obuf/U0/EOUT ));
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_10  (.A(VCC)
        , .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/CCC_0/CCC_INST/PLL_ARST_N_net ), .IPB(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX2_HOLD_N_net ), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_209  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_6  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\demo_sb_sb_0/CCC_0/CCC_INST/CLK2_net ), 
        .IPB(), .IPC(\demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[4] ));
    IOBI_IB_OB_EB \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD/U_IOBI  
        (.D(VCC), .E(VCC), .YIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_126  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] )
        , .IPC());
    IOOUTFF_BYPASS \BIBUF_0/U0/U_IOOUTFF  (.A(\BIBUF_0/U0/DOUT1 ), .Y(
        \BIBUF_0/U0/DOUT ));
    IOBI_IB_OB_EB \BIBUF_0/U0/U_IOBI  (.D(demo_sb_sb_0_I2C_0_SDA_M2F), 
        .E(demo_sb_sb_0_I2C_0_SDA_M2F_OE), .YIN(\BIBUF_0/U0/YIN ), 
        .DOUT(\BIBUF_0/U0/DOUT1 ), .EOUT(\BIBUF_0/U0/EOUT1 ), .Y(
        BIBUF_0_Y));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_252  
        (.A(VCC), .B(VCC), .C(GND), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_16  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_36  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_10  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_30  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_163  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_7  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\demo_sb_sb_0/CCC_0/CCC_INST/CLK3_net ), 
        .IPB(), .IPC(\demo_sb_sb_0/CCC_0/CCC_INST/PWDATA_net[5] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_254  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] )
        , .IPC());
    IOENFF_BYPASS \GPIO_3_M2F_obuf/U0/U_IOENFF  (.A(
        \GPIO_3_M2F_obuf/U0/EOUT1 ), .Y(\GPIO_3_M2F_obuf/U0/EOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_103  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[3] ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net ), 
        .IPC());
    IOOUTFF_BYPASS \GPIO_8_M2F_obuf/U0/U_IOOUTFF  (.A(
        \GPIO_8_M2F_obuf/U0/DOUT1 ), .Y(\GPIO_8_M2F_obuf/U0/DOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_216  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_255  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_83  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_26  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_282  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_84  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[0] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_20  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net )
        , .IPC());
    IOTRI_OB_EB \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DO_PAD/U_IOOUT  (
        .D(VCC), .E(VCC), .DOUT(), .EOUT());
    IOTRI_OB_EB \GPIO_8_M2F_obuf/U0/U_IOTRI  (.D(GPIO_8_M2F_c), .E(VCC)
        , .DOUT(\GPIO_8_M2F_obuf/U0/DOUT1 ), .EOUT(
        \GPIO_8_M2F_obuf/U0/EOUT1 ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_61  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_55  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_284  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] )
        , .IPC());
    IOOUTFF_BYPASS \GPIO_3_M2F_obuf/U0/U_IOOUTFF  (.A(
        \GPIO_3_M2F_obuf/U0/DOUT1 ), .Y(\GPIO_3_M2F_obuf/U0/DOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_178  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net )
        , .IPC());
    SLE \demo_sb_sb_0/CORERESETP_0/RESET_N_F2M_int  (.D(VCC), .CLK(
        \demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1 ), .EN(
        VCC), .ALn(
        \demo_sb_sb_0/CORERESETP_0/POWER_ON_RESET_N_clk_base_Z ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \demo_sb_sb_0/CORERESETP_0_RESET_N_F2M ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_162  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_135  
        (.A(VCC), .B(\demo_sb_sb_0/CORERESETP_0_RESET_N_F2M ), .C(VCC), 
        .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net )
        , .IPC());
    IOBI_IB_OB_EB \BIBUF_1/U0/U_IOBI  (.D(demo_sb_sb_0_I2C_0_SCL_M2F), 
        .E(demo_sb_sb_0_I2C_0_SCL_M2F_OE), .YIN(\BIBUF_1/U0/YIN ), 
        .DOUT(\BIBUF_1/U0/DOUT1 ), .EOUT(\BIBUF_1/U0/EOUT1 ), .Y(
        BIBUF_1_Y));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_145  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_102  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[2] ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[9] ), 
        .IPC());
    GBM_NG \demo_sb_sb_0/CCC_0/GL0_INST  (.An(AFLSDF_INV_0_net_1), 
        .ENn(GND), .YWn(), .YEn(
        \demo_sb_sb_0/CCC_0/GL0_INST/U0_YWn_GEast ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_277  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_116  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_99  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[6] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_59  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_285  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_137  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] )
        , .IPC());
    IP_INTERFACE \demo_sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_12  (.A(VCC)
        , .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/CCC_0/CCC_INST/NGMUX0_ARST_N_net ), .IPB(), .IPC(
        \demo_sb_sb_0/CCC_0/CCC_INST/PADDR_net[2] ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_279  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_147  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_128  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_98  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDIF_net ), .IPB(
        ), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_58  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] )
        , .IPC());
    RGB_NG \demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0  (.An(
        \demo_sb_sb_0/CCC_0/GL0_INST/U0_YWn_GEast ), .ENn(GND), .YL(), 
        .YR(\demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1 ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_17  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_37  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_227  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] )
        , .IPC());
    IOBI_IB_OB_EB \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD/U_IOBI  
        (.D(VCC), .E(VCC), .YIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_263  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_229  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_173  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_203  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_169  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_161  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_109  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_101  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[1] ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[8] ), 
        .IPC());
    SLE \demo_sb_sb_0/CORERESETP_0/POWER_ON_RESET_N_clk_base  (.D(
        \demo_sb_sb_0/CORERESETP_0/sm1_areset_n_q1_Z ), .CLK(
        \demo_sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1 ), .EN(
        VCC), .ALn(\demo_sb_sb_0/SYSRESET_POR_Z ), .ADn(VCC), .SLn(VCC)
        , .SD(GND), .LAT(GND), .Q(
        \demo_sb_sb_0/CORERESETP_0/POWER_ON_RESET_N_clk_base_Z ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_164  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_12  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_32  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_261  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_104  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[4] ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_27  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_201  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_123  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_238  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_248  
        (.A(VCC), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_160  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net )
        , .IPC());
    IOTRI_OB_EB \MMUART_0_TXD_M2F_obuf/U0/U_IOTRI  (.D(
        MMUART_0_TXD_M2F_c), .E(VCC), .DOUT(
        \MMUART_0_TXD_M2F_obuf/U0/DOUT1 ), .EOUT(
        \MMUART_0_TXD_M2F_obuf/U0/EOUT1 ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_100  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[0] ), 
        .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[7] ), 
        .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_45  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_172  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_22  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] )
        , .IPC());
    MSS_025_IP #( .INIT(1438'h0000300C000000300000000000000000000000000000000000000000000000000000000000000000000000000000000001203610000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33F00000000E094C0700003FFFFE4000000000000100000000F0F01C000001825D44010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.000000), .RTC_MAIN_XTL_MODE(""), .DDR_CLK_FREQ(100.000000)
         )  
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/INST_MSS_025_IP  
        (.CAN_RXBUS_MGPIO3A_H2F_A(), .CAN_RXBUS_MGPIO3A_H2F_B(
        GPIO_3_M2F_c), .CAN_TX_EBL_MGPIO4A_H2F_A(), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(GPIO_4_M2F_c), 
        .CAN_TXBUS_MGPIO2A_H2F_A(), .CAN_TXBUS_MGPIO2A_H2F_B(
        GPIO_2_M2F_c), .CLK_CONFIG_APB(), .COMMS_INT(), 
        .CONFIG_PRESET_N(), .EDAC_ERROR({nc16, nc17, nc18, nc19, nc20, 
        nc21, nc22, nc23}), .F_FM0_RDATA({nc24, nc25, nc26, nc27, nc28, 
        nc29, nc30, nc31, nc32, nc33, nc34, nc35, nc36, nc37, nc38, 
        nc39, nc40, nc41, nc42, nc43, nc44, nc45, nc46, nc47, nc48, 
        nc49, nc50, nc51, nc52, nc53, nc54, nc55}), .F_FM0_READYOUT(), 
        .F_FM0_RESP(), .F_HM0_ADDR({nc56, nc57, nc58, nc59, nc60, nc61, 
        nc62, nc63, nc64, nc65, nc66, nc67, nc68, nc69, nc70, nc71, 
        nc72, nc73, nc74, nc75, nc76, nc77, nc78, nc79, nc80, nc81, 
        nc82, nc83, nc84, nc85, nc86, nc87}), .F_HM0_ENABLE(), 
        .F_HM0_SEL(), .F_HM0_SIZE({nc88, nc89}), .F_HM0_TRANS1(), 
        .F_HM0_WDATA({nc90, nc91, nc92, nc93, nc94, nc95, nc96, nc97, 
        nc98, nc99, nc100, nc101, nc102, nc103, nc104, nc105, nc106, 
        nc107, nc108, nc109, nc110, nc111, nc112, nc113, nc114, nc115, 
        nc116, nc117, nc118, nc119, nc120, nc121}), .F_HM0_WRITE(), 
        .FAB_CHRGVBUS(), .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), 
        .FAB_DPPULLDOWN(), .FAB_DRVVBUS(), .FAB_IDPULLUP(), 
        .FAB_OPMODE({nc122, nc123}), .FAB_SUSPENDM(), .FAB_TERMSEL(), 
        .FAB_TXVALID(), .FAB_VCONTROL({nc124, nc125, nc126, nc127}), 
        .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({nc128, nc129}), 
        .FAB_XDATAOUT({nc130, nc131, nc132, nc133, nc134, nc135, nc136, 
        nc137}), .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc138, nc139}), 
        .FIC32_1_MASTER({nc140, nc141}), .FPGA_RESET_N(), .GTX_CLK(), 
        .H2F_INTERRUPT({nc142, nc143, nc144, nc145, nc146, nc147, 
        nc148, nc149, nc150, nc151, nc152, nc153, nc154, nc155, nc156, 
        nc157}), .H2F_NMI(), .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(
        demo_sb_sb_0_I2C_0_SCL_M2F), .I2C0_SCL_MGPIO31B_H2F_B(
        demo_sb_sb_0_I2C_0_SCL_M2F_OE), .I2C0_SDA_MGPIO30B_H2F_A(
        demo_sb_sb_0_I2C_0_SDA_M2F), .I2C0_SDA_MGPIO30B_H2F_B(
        demo_sb_sb_0_I2C_0_SDA_M2F_OE), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(), .I2C1_SDA_MGPIO0A_H2F_A(), 
        .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), .MDOENF(), .MDOF(), 
        .MMUART0_CTS_MGPIO19B_H2F_A(), .MMUART0_CTS_MGPIO19B_H2F_B(), 
        .MMUART0_DCD_MGPIO22B_H2F_A(), .MMUART0_DCD_MGPIO22B_H2F_B(), 
        .MMUART0_DSR_MGPIO20B_H2F_A(), .MMUART0_DSR_MGPIO20B_H2F_B(), 
        .MMUART0_DTR_MGPIO18B_H2F_A(), .MMUART0_DTR_MGPIO18B_H2F_B(), 
        .MMUART0_RI_MGPIO21B_H2F_A(), .MMUART0_RI_MGPIO21B_H2F_B(), 
        .MMUART0_RTS_MGPIO17B_H2F_A(), .MMUART0_RTS_MGPIO17B_H2F_B(), 
        .MMUART0_RXD_MGPIO28B_H2F_A(), .MMUART0_RXD_MGPIO28B_H2F_B(), 
        .MMUART0_SCK_MGPIO29B_H2F_A(), .MMUART0_SCK_MGPIO29B_H2F_B(), 
        .MMUART0_TXD_MGPIO27B_H2F_A(MMUART_0_TXD_M2F_c), 
        .MMUART0_TXD_MGPIO27B_H2F_B(), .MMUART1_DTR_MGPIO12B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_B(), 
        .MMUART1_RXD_MGPIO26B_H2F_A(), .MMUART1_RXD_MGPIO26B_H2F_B(), 
        .MMUART1_SCK_MGPIO25B_H2F_A(), .MMUART1_SCK_MGPIO25B_H2F_B(), 
        .MMUART1_TXD_MGPIO24B_H2F_A(), .MMUART1_TXD_MGPIO24B_H2F_B(), 
        .MPLL_LOCK(), .PER2_FABRIC_PADDR({nc158, nc159, nc160, nc161, 
        nc162, nc163, nc164, nc165, nc166, nc167, nc168, nc169, nc170, 
        nc171}), .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc172, nc173, nc174, nc175, nc176, nc177, 
        nc178, nc179, nc180, nc181, nc182, nc183, nc184, nc185, nc186, 
        nc187, nc188, nc189, nc190, nc191, nc192, nc193, nc194, nc195, 
        nc196, nc197, nc198, nc199, nc200, nc201, nc202, nc203}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(
        GPIO_8_M2F_c), .SPI0_SS2_MGPIO9A_H2F_A(), 
        .SPI0_SS2_MGPIO9A_H2F_B(), .SPI0_SS3_MGPIO10A_H2F_A(), 
        .SPI0_SS3_MGPIO10A_H2F_B(), .SPI0_SS4_MGPIO19A_H2F_A(), 
        .SPI0_SS5_MGPIO20A_H2F_A(), .SPI0_SS6_MGPIO21A_H2F_A(), 
        .SPI0_SS7_MGPIO22A_H2F_A(), .SPI1_CLK_OUT(), 
        .SPI1_SDI_MGPIO11A_H2F_A(), .SPI1_SDI_MGPIO11A_H2F_B(), 
        .SPI1_SDO_MGPIO12A_H2F_A(), .SPI1_SDO_MGPIO12A_H2F_B(), 
        .SPI1_SS0_MGPIO13A_H2F_A(), .SPI1_SS0_MGPIO13A_H2F_B(), 
        .SPI1_SS1_MGPIO14A_H2F_A(), .SPI1_SS1_MGPIO14A_H2F_B(), 
        .SPI1_SS2_MGPIO15A_H2F_A(), .SPI1_SS2_MGPIO15A_H2F_B(), 
        .SPI1_SS3_MGPIO16A_H2F_A(), .SPI1_SS3_MGPIO16A_H2F_B(), 
        .SPI1_SS4_MGPIO17A_H2F_A(), .SPI1_SS5_MGPIO18A_H2F_A(), 
        .SPI1_SS6_MGPIO23A_H2F_A(), .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({
        nc204, nc205, nc206, nc207, nc208, nc209, nc210, nc211, nc212, 
        nc213}), .TRACECLK(), .TRACEDATA({nc214, nc215, nc216, nc217}), 
        .TX_CLK(), .TX_ENF(), .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({
        nc218, nc219, nc220, nc221}), .TXDF({nc222, nc223, nc224, 
        nc225, nc226, nc227, nc228, nc229}), .TXEV(), .WDOGTIMEOUT(), 
        .F_ARREADY_HREADYOUT1(), .F_AWREADY_HREADYOUT0(), .F_BID({
        nc230, nc231, nc232, nc233}), .F_BRESP_HRESP0({nc234, nc235}), 
        .F_BVALID(), .F_RDATA_HRDATA01({nc236, nc237, nc238, nc239, 
        nc240, nc241, nc242, nc243, nc244, nc245, nc246, nc247, nc248, 
        nc249, nc250, nc251, nc252, nc253, nc254, nc255, nc256, nc257, 
        nc258, nc259, nc260, nc261, nc262, nc263, nc264, nc265, nc266, 
        nc267, nc268, nc269, nc270, nc271, nc272, nc273, nc274, nc275, 
        nc276, nc277, nc278, nc279, nc280, nc281, nc282, nc283, nc284, 
        nc285, nc286, nc287, nc288, nc289, nc290, nc291, nc292, nc293, 
        nc294, nc295, nc296, nc297, nc298, nc299}), .F_RID({nc300, 
        nc301, nc302, nc303}), .F_RLAST(), .F_RRESP_HRESP1({nc304, 
        nc305}), .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc306, 
        nc307, nc308, nc309, nc310, nc311, nc312, nc313, nc314, nc315, 
        nc316, nc317, nc318, nc319, nc320, nc321}), 
        .MDDR_FABRIC_PREADY(), .MDDR_FABRIC_PSLVERR(), 
        .CAN_RXBUS_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net )
        , .CAN_TX_EBL_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net )
        , .CAN_TXBUS_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net )
        , .COLF(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/COLF_net ), 
        .CRSF(\demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CRSF_net ), 
        .F2_DMAREADY({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] })
        , .F2H_INTERRUPT({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] })
        , .F2HCALIB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F2HCALIB_net ), 
        .F_DMAREADY({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] })
        , .F_FM0_ADDR({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] })
        , .F_FM0_ENABLE(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net )
        , .F_FM0_MASTLOCK(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net )
        , .F_FM0_READY(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net )
        , .F_FM0_SEL(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net ), 
        .F_FM0_SIZE({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] })
        , .F_FM0_TRANS1(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net )
        , .F_FM0_WDATA({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] })
        , .F_FM0_WRITE(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net )
        , .F_HM0_RDATA({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] })
        , .F_HM0_READY(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net )
        , .F_HM0_RESP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net ), 
        .FAB_AVALID(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net ), 
        .FAB_HOSTDISCON(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net )
        , .FAB_IDDIG(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net ), 
        .FAB_LINESTATE({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] })
        , .FAB_M3_RESET_N(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net )
        , .FAB_PLL_LOCK(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net )
        , .FAB_RXACTIVE(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net )
        , .FAB_RXERROR(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net )
        , .FAB_RXVALID(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net )
        , .FAB_RXVALIDH(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net )
        , .FAB_SESSEND(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net )
        , .FAB_TXREADY(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net )
        , .FAB_VBUSVALID(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net )
        , .FAB_VSTATUS({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] })
        , .FAB_XDATAIN({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] })
        , .GTX_CLKPF(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net ), 
        .I2C0_BCLK(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net ), 
        .I2C0_SCL_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net )
        , .I2C0_SDA_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net )
        , .I2C1_BCLK(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net ), 
        .I2C1_SCL_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net )
        , .I2C1_SDA_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net )
        , .MDIF(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDIF_net ), 
        .MGPIO0A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net )
        , .MGPIO10A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net )
        , .MGPIO11A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net )
        , .MGPIO11B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net )
        , .MGPIO12A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net )
        , .MGPIO13A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net )
        , .MGPIO14A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net )
        , .MGPIO15A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net )
        , .MGPIO16A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net )
        , .MGPIO17B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net )
        , .MGPIO18B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net )
        , .MGPIO19B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net )
        , .MGPIO1A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net )
        , .MGPIO20B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net )
        , .MGPIO21B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net )
        , .MGPIO22B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net )
        , .MGPIO24B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net )
        , .MGPIO25B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net )
        , .MGPIO26B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net )
        , .MGPIO27B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net )
        , .MGPIO28B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net )
        , .MGPIO29B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net )
        , .MGPIO2A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net )
        , .MGPIO30B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net )
        , .MGPIO31B_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net )
        , .MGPIO3A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net )
        , .MGPIO4A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net )
        , .MGPIO5A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net )
        , .MGPIO6A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net )
        , .MGPIO7A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net )
        , .MGPIO8A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net )
        , .MGPIO9A_F2H_GPIN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net )
        , .MMUART0_CTS_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net )
        , .MMUART0_DCD_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net )
        , .MMUART0_DSR_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net )
        , .MMUART0_DTR_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net )
        , .MMUART0_RI_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net )
        , .MMUART0_RTS_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net )
        , .MMUART0_RXD_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net )
        , .MMUART0_SCK_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net )
        , .MMUART0_TXD_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net )
        , .MMUART1_CTS_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net )
        , .MMUART1_DCD_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net )
        , .MMUART1_DSR_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net )
        , .MMUART1_RI_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net )
        , .MMUART1_RTS_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net )
        , .MMUART1_RXD_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net )
        , .MMUART1_SCK_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net )
        , .MMUART1_TXD_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net )
        , .PER2_FABRIC_PRDATA({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] })
        , .PER2_FABRIC_PREADY(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net )
        , .PER2_FABRIC_PSLVERR(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net )
        , .RCGF({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[0] }), 
        .RX_CLKPF(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net ), 
        .RX_DVF(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_DVF_net ), 
        .RX_ERRF(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_ERRF_net ), 
        .RX_EV(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RX_EV_net ), 
        .RXDF({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[0] }), 
        .SLEEPHOLDREQ(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net )
        , .SMBALERT_NI0(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net )
        , .SMBALERT_NI1(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net )
        , .SMBSUS_NI0(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net ), 
        .SMBSUS_NI1(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net ), 
        .SPI0_CLK_IN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net )
        , .SPI0_SDI_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net )
        , .SPI0_SDO_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net )
        , .SPI0_SS0_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net )
        , .SPI0_SS1_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net )
        , .SPI0_SS2_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net )
        , .SPI0_SS3_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net )
        , .SPI1_CLK_IN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net )
        , .SPI1_SDI_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net )
        , .SPI1_SDO_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net )
        , .SPI1_SS0_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net )
        , .SPI1_SS1_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net )
        , .SPI1_SS2_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net )
        , .SPI1_SS3_F2H_SCP(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net )
        , .TX_CLKPF(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net ), 
        .USER_MSS_GPIO_RESET_N(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net )
        , .USER_MSS_RESET_N(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net )
        , .XCLK_FAB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net ), 
        .CLK_BASE(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CLK_BASE_net ), 
        .CLK_MDDR_APB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net )
        , .F_ARADDR_HADDR1({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] })
        , .F_ARBURST_HTRANS1({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] })
        , .F_ARID_HSEL1({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] })
        , .F_ARLEN_HBURST1({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] })
        , .F_ARLOCK_HMASTLOCK1({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] })
        , .F_ARSIZE_HSIZE1({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] })
        , .F_ARVALID_HWRITE1(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net )
        , .F_AWADDR_HADDR0({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] })
        , .F_AWBURST_HTRANS0({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] })
        , .F_AWID_HSEL0({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] })
        , .F_AWLEN_HBURST0({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] })
        , .F_AWLOCK_HMASTLOCK0({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] })
        , .F_AWSIZE_HSIZE0({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] })
        , .F_AWVALID_HWRITE0(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net )
        , .F_BREADY(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_BREADY_net ), 
        .F_RMW_AXI(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net ), 
        .F_RREADY(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_RREADY_net ), 
        .F_WDATA_HWDATA01({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] })
        , .F_WID_HREADY01({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] })
        , .F_WLAST(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WLAST_net ), 
        .F_WSTRB({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] })
        , .F_WVALID(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WVALID_net ), 
        .FPGA_MDDR_ARESET_N(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net )
        , .MDDR_FABRIC_PADDR({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] })
        , .MDDR_FABRIC_PENABLE(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net )
        , .MDDR_FABRIC_PSEL(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net )
        , .MDDR_FABRIC_PWDATA({
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] , 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] })
        , .MDDR_FABRIC_PWRITE(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net )
        , .PRESET_N(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PRESET_N_net ), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND), .DM_IN({GND, GND, GND}), 
        .DRAM_DQ_IN({GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .DRAM_DQS_IN({GND, 
        GND, GND}), .DRAM_FIFO_WE_IN({GND, GND}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND), .MGPIO25A_IN(GND), 
        .MGPIO26A_IN(GND), .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND), 
        .MMUART0_DCD_MGPIO22B_IN(GND), .MMUART0_DSR_MGPIO20B_IN(GND), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND), 
        .MMUART0_RI_MGPIO21B_IN(GND), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(GND), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND), 
        .MMUART1_CTS_MGPIO13B_IN(GND), .MMUART1_DCD_MGPIO16B_IN(GND), 
        .MMUART1_DSR_MGPIO14B_IN(GND), .MMUART1_DTR_MGPIO12B_IN(GND), 
        .MMUART1_RI_MGPIO15B_IN(GND), .MMUART1_RTS_MGPIO11B_IN(GND), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND), 
        .RGMII_MDC_RMII_MDC_IN(GND), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND), .RGMII_RX_CLK_IN(GND)
        , .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND), 
        .RGMII_RXD3_USBB_DATA4_IN(GND), .RGMII_TX_CLK_IN(GND), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND), 
        .RGMII_TXD2_USBB_DATA5_IN(GND), .RGMII_TXD3_USBB_DATA6_IN(GND), 
        .SPI0_SCK_USBA_XCLK_IN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD_Y ), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_IN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DI_PAD_Y ), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_SS0_PAD_Y ), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND), .SPI0_SS4_MGPIO19A_IN(
        GND), .SPI0_SS5_MGPIO20A_IN(GND), .SPI0_SS6_MGPIO21A_IN(GND), 
        .SPI0_SS7_MGPIO22A_IN(GND), .SPI1_SCK_IN(GND), 
        .SPI1_SDI_MGPIO11A_IN(GND), .SPI1_SDO_MGPIO12A_IN(GND), 
        .SPI1_SS0_MGPIO13A_IN(GND), .SPI1_SS1_MGPIO14A_IN(GND), 
        .SPI1_SS2_MGPIO15A_IN(GND), .SPI1_SS3_MGPIO16A_IN(GND), 
        .SPI1_SS4_MGPIO17A_IN(GND), .SPI1_SS5_MGPIO18A_IN(GND), 
        .SPI1_SS6_MGPIO23A_IN(GND), .SPI1_SS7_MGPIO24A_IN(GND), 
        .USBC_XCLK_IN(GND), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc322, nc323, 
        nc324, nc325, nc326, nc327, nc328, nc329, nc330, nc331, nc332, 
        nc333, nc334, nc335, nc336, nc337}), .DRAM_BA({nc338, nc339, 
        nc340}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc341, nc342, nc343}), .DRAM_DQ_OUT({nc344, 
        nc345, nc346, nc347, nc348, nc349, nc350, nc351, nc352, nc353, 
        nc354, nc355, nc356, nc357, nc358, nc359, nc360, nc361}), 
        .DRAM_DQS_OUT({nc362, nc363, nc364}), .DRAM_FIFO_WE_OUT({nc365, 
        nc366}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), .MGPIO25A_OUT(), 
        .MGPIO26A_OUT(), .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(), 
        .MMUART1_CTS_MGPIO13B_OUT(), .MMUART1_DCD_MGPIO16B_OUT(), 
        .MMUART1_DSR_MGPIO14B_OUT(), .MMUART1_DTR_MGPIO12B_OUT(), 
        .MMUART1_RI_MGPIO15B_OUT(), .MMUART1_RTS_MGPIO11B_OUT(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT )
        , .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT )
        , .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT )
        , .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI0_SS4_MGPIO19A_OUT(), 
        .SPI0_SS5_MGPIO20A_OUT(), .SPI0_SS6_MGPIO21A_OUT(), 
        .SPI0_SS7_MGPIO22A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc367, nc368, 
        nc369}), .DRAM_DQ_OE({nc370, nc371, nc372, nc373, nc374, nc375, 
        nc376, nc377, nc378, nc379, nc380, nc381, nc382, nc383, nc384, 
        nc385, nc386, nc387}), .DRAM_DQS_OE({nc388, nc389, nc390}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), .MGPIO25A_OE(), 
        .MGPIO26A_OE(), .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(), .MMUART1_CTS_MGPIO13B_OE()
        , .MMUART1_DCD_MGPIO16B_OE(), .MMUART1_DSR_MGPIO14B_OE(), 
        .MMUART1_DTR_MGPIO12B_OE(), .MMUART1_RI_MGPIO15B_OE(), 
        .MMUART1_RTS_MGPIO11B_OE(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE )
        , .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE )
        , .SPI0_SS0_USBA_NXT_MGPIO7A_OE(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE )
        , .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI0_SS4_MGPIO19A_OE(), 
        .SPI0_SS5_MGPIO20A_OE(), .SPI0_SS6_MGPIO21A_OE(), 
        .SPI0_SS7_MGPIO22A_OE(), .SPI1_SCK_OE(), .SPI1_SDI_MGPIO11A_OE(
        ), .SPI1_SDO_MGPIO12A_OE(), .SPI1_SS0_MGPIO13A_OE(), 
        .SPI1_SS1_MGPIO14A_OE(), .SPI1_SS2_MGPIO15A_OE(), 
        .SPI1_SS3_MGPIO16A_OE(), .SPI1_SS4_MGPIO17A_OE(), 
        .SPI1_SS5_MGPIO18A_OE(), .SPI1_SS6_MGPIO23A_OE(), 
        .SPI1_SS7_MGPIO24A_OE(), .USBC_XCLK_OE());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_6  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_118  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_75  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_230  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_49  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_217  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] )
        , .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_240  
        (.A(VCC), .B(GND), .C(GND), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] ), 
        .IPC(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WVALID_net ));
    IOENFF_BYPASS \GPIO_8_M2F_obuf/U0/U_IOENFF  (.A(
        \GPIO_8_M2F_obuf/U0/EOUT1 ), .Y(\GPIO_8_M2F_obuf/U0/EOUT ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_219  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] )
        , .IPC());
    sdf_IOPAD_BI \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD/U_IOPAD  
        (.PAD(SPI_0_CLK), .D(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT )
        , .E(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE )
        , .Y(\demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_CLK_PAD_Y ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_122  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net )
        , .IPB(), .IPC());
    IOTRI_OB_EB \GPIO_2_M2F_obuf/U0/U_IOTRI  (.D(GPIO_2_M2F_c), .E(VCC)
        , .DOUT(\GPIO_2_M2F_obuf/U0/DOUT1 ), .EOUT(
        \GPIO_2_M2F_obuf/U0/EOUT1 ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_79  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_48  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] )
        , .IPB(), .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_273  
        (.A(GND), .B(VCC), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net )
        , .IPC());
    IOTRI_OB_EB \GPIO_4_M2F_obuf/U0/U_IOTRI  (.D(GPIO_4_M2F_c), .E(VCC)
        , .DOUT(\GPIO_4_M2F_obuf/U0/DOUT1 ), .EOUT(
        \GPIO_4_M2F_obuf/U0/EOUT1 ));
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_11  
        (.A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] )
        , .IPC());
    sdf_IOPAD_TRI \demo_sb_sb_0/demo_sb_sb_MSS_0/SPI_0_DO_PAD/U_IOPAD  
        (.PAD(SPI_0_DO), .D(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT )
        , .E(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE )
        );
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_31  
        (.A(GND), .B(GND), .C(VCC), .IPA(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] )
        , .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] )
        , .IPC());
    IP_INTERFACE 
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_179  
        (.A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \demo_sb_sb_0/demo_sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net )
        , .IPC());
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
